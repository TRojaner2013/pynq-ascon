// Message Types for communicaton with PS.
`define KEY 4'd0
`define NONCE 4'd1
`define AD 4'd2
`define PLAIN 4'd3
`define CIPHER 4'd4
`define TAG 4'd5
`define MSG 4'd6
`define HASH 4'd7
`define LEN 4'd8
`define CONF 4'd9
`define ABORT 4'd10
`define OK 4'd11
`define SKIP_AD 4'd12
